mem[0] = "\033";
mem[1] = "[";
mem[2] = "2";
mem[3] = "J";
mem[4] = "\033";
mem[5] = "[";
mem[6] = "1";
mem[7] = ";";
mem[8] = "1";
mem[9] = "H";
mem[10] = "\015";
mem[11] = "\012";
mem[12] = "R";
mem[13] = "e";
mem[14] = "a";
mem[15] = "d";
mem[16] = "y";
mem[17] = "\015";
mem[18] = "\012";
mem[19] = "\033";
mem[20] = "[";
mem[21] = "0";
mem[22] = "2";
mem[23] = "m";
mem[24] = " ";
mem[25] = " ";
mem[26] = " ";
mem[27] = " ";
mem[28] = " ";
mem[29] = " ";
mem[30] = "t";
mem[31] = "x";
mem[32] = "_";
mem[33] = "e";
mem[34] = "n";
mem[35] = " ";
mem[36] = " ";
mem[37] = " ";
mem[38] = " ";
mem[39] = " ";
mem[40] = " ";
mem[41] = " ";
mem[42] = " ";
mem[43] = " ";
mem[44] = "\033";
mem[45] = "[";
mem[46] = "0";
mem[47] = "0";
mem[48] = "m";
mem[49] = "\015";
mem[50] = "\012";
mem[51] = "\033";
mem[52] = "[";
mem[53] = "0";
mem[54] = "2";
mem[55] = "m";
mem[56] = " ";
mem[57] = " ";
mem[58] = " ";
mem[59] = " ";
mem[60] = " ";
mem[61] = " ";
mem[62] = " ";
mem[63] = "t";
mem[64] = "x";
mem[65] = "_";
mem[66] = "j";
mem[67] = " ";
mem[68] = " ";
mem[69] = " ";
mem[70] = " ";
mem[71] = " ";
mem[72] = " ";
mem[73] = " ";
mem[74] = " ";
mem[75] = " ";
mem[76] = "\033";
mem[77] = "[";
mem[78] = "0";
mem[79] = "0";
mem[80] = "m";
mem[81] = "\015";
mem[82] = "\012";
mem[83] = "\033";
mem[84] = "[";
mem[85] = "0";
mem[86] = "2";
mem[87] = "m";
mem[88] = " ";
mem[89] = " ";
mem[90] = " ";
mem[91] = " ";
mem[92] = " ";
mem[93] = " ";
mem[94] = "t";
mem[95] = "x";
mem[96] = "_";
mem[97] = "s";
mem[98] = "e";
mem[99] = "0";
mem[100] = " ";
mem[101] = " ";
mem[102] = " ";
mem[103] = " ";
mem[104] = " ";
mem[105] = " ";
mem[106] = " ";
mem[107] = " ";
mem[108] = "\033";
mem[109] = "[";
mem[110] = "0";
mem[111] = "0";
mem[112] = "m";
mem[113] = "\015";
mem[114] = "\012";
mem[115] = "\033";
mem[116] = "[";
mem[117] = "0";
mem[118] = "2";
mem[119] = "m";
mem[120] = " ";
mem[121] = " ";
mem[122] = " ";
mem[123] = " ";
mem[124] = " ";
mem[125] = " ";
mem[126] = "u";
mem[127] = "s";
mem[128] = "b";
mem[129] = "_";
mem[130] = "r";
mem[131] = "s";
mem[132] = "t";
mem[133] = " ";
mem[134] = " ";
mem[135] = " ";
mem[136] = " ";
mem[137] = " ";
mem[138] = " ";
mem[139] = " ";
mem[140] = "\033";
mem[141] = "[";
mem[142] = "0";
mem[143] = "0";
mem[144] = "m";
mem[145] = "\015";
mem[146] = "\012";
mem[147] = "\033";
mem[148] = "[";
mem[149] = "0";
mem[150] = "2";
mem[151] = "m";
mem[152] = " ";
mem[153] = "t";
mem[154] = "r";
mem[155] = "a";
mem[156] = "n";
mem[157] = "s";
mem[158] = "a";
mem[159] = "c";
mem[160] = "t";
mem[161] = "i";
mem[162] = "o";
mem[163] = "n";
mem[164] = "_";
mem[165] = "a";
mem[166] = "c";
mem[167] = "t";
mem[168] = "i";
mem[169] = "v";
mem[170] = "e";
mem[171] = " ";
mem[172] = "\033";
mem[173] = "[";
mem[174] = "0";
mem[175] = "0";
mem[176] = "m";
mem[177] = "\015";
mem[178] = "\012";
mem[179] = "\033";
mem[180] = "[";
mem[181] = "0";
mem[182] = "0";
mem[183] = "m";
mem[184] = " ";
mem[185] = " ";
mem[186] = " ";
mem[187] = " ";
mem[188] = " ";
mem[189] = "e";
mem[190] = "n";
mem[191] = "d";
mem[192] = "p";
mem[193] = "o";
mem[194] = "i";
mem[195] = "n";
mem[196] = "t";
mem[197] = ":";
mem[198] = " ";
mem[199] = "0";
mem[200] = " ";
mem[201] = " ";
mem[202] = " ";
mem[203] = " ";
mem[204] = "\033";
mem[205] = "[";
mem[206] = "0";
mem[207] = "0";
mem[208] = "m";
mem[209] = "\015";
mem[210] = "\012";
mem[211] = "\033";
mem[212] = "[";
mem[213] = "0";
mem[214] = "2";
mem[215] = "m";
mem[216] = " ";
mem[217] = " ";
mem[218] = " ";
mem[219] = " ";
mem[220] = "d";
mem[221] = "i";
mem[222] = "r";
mem[223] = "e";
mem[224] = "c";
mem[225] = "t";
mem[226] = "i";
mem[227] = "o";
mem[228] = "n";
mem[229] = "_";
mem[230] = "i";
mem[231] = "n";
mem[232] = " ";
mem[233] = " ";
mem[234] = " ";
mem[235] = " ";
mem[236] = "\033";
mem[237] = "[";
mem[238] = "0";
mem[239] = "0";
mem[240] = "m";
mem[241] = "\015";
mem[242] = "\012";
mem[243] = "\033";
mem[244] = "[";
mem[245] = "0";
mem[246] = "2";
mem[247] = "m";
mem[248] = " ";
mem[249] = " ";
mem[250] = " ";
mem[251] = " ";
mem[252] = " ";
mem[253] = " ";
mem[254] = " ";
mem[255] = "s";
mem[256] = "e";
mem[257] = "t";
mem[258] = "u";
mem[259] = "p";
mem[260] = " ";
mem[261] = " ";
mem[262] = " ";
mem[263] = " ";
mem[264] = " ";
mem[265] = " ";
mem[266] = " ";
mem[267] = " ";
mem[268] = "\033";
mem[269] = "[";
mem[270] = "0";
mem[271] = "0";
mem[272] = "m";
mem[273] = "\015";
mem[274] = "\012";
mem[275] = "\033";
mem[276] = "[";
mem[277] = "0";
mem[278] = "2";
mem[279] = "m";
mem[280] = " ";
mem[281] = " ";
mem[282] = " ";
mem[283] = " ";
mem[284] = "d";
mem[285] = "a";
mem[286] = "t";
mem[287] = "a";
mem[288] = "_";
mem[289] = "s";
mem[290] = "t";
mem[291] = "r";
mem[292] = "o";
mem[293] = "b";
mem[294] = "e";
mem[295] = " ";
mem[296] = " ";
mem[297] = " ";
mem[298] = " ";
mem[299] = " ";
mem[300] = "\033";
mem[301] = "[";
mem[302] = "0";
mem[303] = "0";
mem[304] = "m";
mem[305] = "\015";
mem[306] = "\012";
mem[307] = "\033";
mem[308] = "[";
mem[309] = "0";
mem[310] = "2";
mem[311] = "m";
mem[312] = " ";
mem[313] = " ";
mem[314] = " ";
mem[315] = " ";
mem[316] = " ";
mem[317] = " ";
mem[318] = "s";
mem[319] = "u";
mem[320] = "c";
mem[321] = "c";
mem[322] = "e";
mem[323] = "s";
mem[324] = "s";
mem[325] = " ";
mem[326] = " ";
mem[327] = " ";
mem[328] = " ";
mem[329] = " ";
mem[330] = " ";
mem[331] = " ";
mem[332] = "\033";
mem[333] = "[";
mem[334] = "0";
mem[335] = "0";
mem[336] = "m";
mem[337] = "\015";
mem[338] = "\012";
mem[339] = "\015";
mem[340] = "\012";
mem[341] = "d";
mem[342] = "a";
mem[343] = "t";
mem[344] = "a";
mem[345] = ":";
mem[346] = "\015";
mem[347] = "\012";
