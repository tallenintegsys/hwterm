mem[0] = " ";
mem[1] = " ";
mem[2] = " ";
mem[3] = " ";
mem[4] = " ";
mem[5] = " ";
mem[6] = " ";
mem[7] = " ";
mem[8] = " ";
mem[9] = " ";
mem[10] = " ";
mem[11] = " ";
mem[12] = " ";
mem[13] = " ";
mem[14] = " ";
mem[15] = " ";
mem[16] = " ";
mem[17] = " ";
mem[18] = " ";
mem[19] = " ";
mem[20] = " ";
mem[21] = "_";
mem[22] = "_";
mem[23] = "_";
mem[24] = "_";
mem[25] = "_";
mem[26] = "_";
mem[27] = "_";
mem[28] = "_";
mem[29] = "_";
mem[30] = "_";
mem[31] = "_";
mem[32] = "_";
mem[33] = "_";
mem[34] = "_";
mem[35] = "_";
mem[36] = "_";
mem[37] = " ";
mem[38] = " ";
mem[39] = " ";
mem[40] = "\015";
mem[41] = "\012";
mem[42] = " ";
mem[43] = " ";
mem[44] = " ";
mem[45] = " ";
mem[46] = " ";
mem[47] = " ";
mem[48] = " ";
mem[49] = " ";
mem[50] = " ";
mem[51] = " ";
mem[52] = " ";
mem[53] = " ";
mem[54] = " ";
mem[55] = " ";
mem[56] = " ";
mem[57] = " ";
mem[58] = " ";
mem[59] = " ";
mem[60] = " ";
mem[61] = " ";
mem[62] = "|";
mem[63] = " ";
mem[64] = " ";
mem[65] = " ";
mem[66] = " ";
mem[67] = " ";
mem[68] = " ";
mem[69] = " ";
mem[70] = " ";
mem[71] = " ";
mem[72] = " ";
mem[73] = " ";
mem[74] = " ";
mem[75] = " ";
mem[76] = " ";
mem[77] = " ";
mem[78] = " ";
mem[79] = "|";
mem[80] = " ";
mem[81] = " ";
mem[82] = "\015";
mem[83] = "\012";
mem[84] = " ";
mem[85] = " ";
mem[86] = "d";
mem[87] = "e";
mem[88] = "l";
mem[89] = "a";
mem[90] = "y";
mem[91] = " ";
mem[92] = " ";
mem[93] = "w";
mem[94] = "i";
mem[95] = "d";
mem[96] = "t";
mem[97] = "h";
mem[98] = " ";
mem[99] = " ";
mem[100] = " ";
mem[101] = " ";
mem[102] = " ";
mem[103] = " ";
mem[104] = "|";
mem[105] = " ";
mem[106] = "p";
mem[107] = "u";
mem[108] = "l";
mem[109] = "s";
mem[110] = "e";
mem[111] = " ";
mem[112] = " ";
mem[113] = "w";
mem[114] = "i";
mem[115] = "d";
mem[116] = "t";
mem[117] = "h";
mem[118] = " ";
mem[119] = " ";
mem[120] = " ";
mem[121] = "|";
mem[122] = " ";
mem[123] = " ";
mem[124] = "\015";
mem[125] = "\012";
mem[126] = " ";
mem[127] = " ";
mem[128] = "";
mem[129] = "[";
mem[130] = "1";
mem[131] = "0";
mem[132] = "0";
mem[133] = "m";
mem[134] = " ";
mem[135] = " ";
mem[136] = " ";
mem[137] = " ";
mem[138] = " ";
mem[139] = " ";
mem[140] = " ";
mem[141] = " ";
mem[142] = " ";
mem[143] = " ";
mem[144] = " ";
mem[145] = " ";
mem[146] = "";
mem[147] = "[";
mem[148] = "m";
mem[149] = " ";
mem[150] = "n";
mem[151] = "s";
mem[152] = " ";
mem[153] = " ";
mem[154] = " ";
mem[155] = "|";
mem[156] = " ";
mem[157] = "";
mem[158] = "[";
mem[159] = "1";
mem[160] = "0";
mem[161] = "0";
mem[162] = "m";
mem[163] = " ";
mem[164] = " ";
mem[165] = " ";
mem[166] = " ";
mem[167] = " ";
mem[168] = " ";
mem[169] = " ";
mem[170] = " ";
mem[171] = " ";
mem[172] = " ";
mem[173] = " ";
mem[174] = " ";
mem[175] = "";
mem[176] = "[";
mem[177] = "m";
mem[178] = " ";
mem[179] = "n";
mem[180] = "s";
mem[181] = "|";
mem[182] = " ";
mem[183] = " ";
mem[184] = "\015";
mem[185] = "\012";
mem[186] = "_";
mem[187] = "_";
mem[188] = "_";
mem[189] = "_";
mem[190] = "_";
mem[191] = "_";
mem[192] = "_";
mem[193] = "_";
mem[194] = "_";
mem[195] = "_";
mem[196] = "_";
mem[197] = "_";
mem[198] = "_";
mem[199] = "_";
mem[200] = "_";
mem[201] = "_";
mem[202] = "_";
mem[203] = "_";
mem[204] = "_";
mem[205] = "_";
mem[206] = "|";
mem[207] = " ";
mem[208] = " ";
mem[209] = " ";
mem[210] = " ";
mem[211] = " ";
mem[212] = " ";
mem[213] = " ";
mem[214] = " ";
mem[215] = " ";
mem[216] = " ";
mem[217] = " ";
mem[218] = " ";
mem[219] = " ";
mem[220] = " ";
mem[221] = " ";
mem[222] = " ";
mem[223] = "|";
mem[224] = "_";
mem[225] = "_";
mem[226] = "\015";
mem[227] = "\012";
mem[228] = "\015";
mem[229] = "\012";
mem[230] = " ";
mem[231] = "t";
mem[232] = "a";
mem[233] = "b";
mem[234] = "=";
mem[235] = "f";
mem[236] = "i";
mem[237] = "e";
mem[238] = "l";
mem[239] = "d";
mem[240] = " ";
mem[241] = "s";
mem[242] = "p";
mem[243] = "a";
mem[244] = "c";
mem[245] = "e";
mem[246] = "=";
mem[247] = "r";
mem[248] = "e";
mem[249] = "d";
mem[250] = "r";
mem[251] = "a";
mem[252] = "w";
mem[253] = " ";
mem[254] = "e";
mem[255] = "n";
mem[256] = "t";
mem[257] = "e";
mem[258] = "r";
mem[259] = "=";
mem[260] = "t";
mem[261] = "r";
mem[262] = "i";
mem[263] = "g";
mem[264] = "g";
mem[265] = "e";
mem[266] = "r";
mem[267] = " ";
mem[268] = " ";
mem[269] = " ";
mem[270] = "\015";
mem[271] = "\012";
