mem[0] = "";
mem[1] = "[";
mem[2] = "2";
mem[3] = "J";
mem[4] = " ";
mem[5] = " ";
mem[6] = " ";
mem[7] = " ";
mem[8] = " ";
mem[9] = " ";
mem[10] = " ";
mem[11] = " ";
mem[12] = " ";
mem[13] = " ";
mem[14] = " ";
mem[15] = " ";
mem[16] = " ";
mem[17] = " ";
mem[18] = " ";
mem[19] = " ";
mem[20] = " ";
mem[21] = " ";
mem[22] = " ";
mem[23] = " ";
mem[24] = " ";
mem[25] = " ";
mem[26] = " ";
mem[27] = " ";
mem[28] = " ";
mem[29] = "_";
mem[30] = "_";
mem[31] = "_";
mem[32] = "_";
mem[33] = "_";
mem[34] = "_";
mem[35] = "_";
mem[36] = "_";
mem[37] = "_";
mem[38] = "_";
mem[39] = "_";
mem[40] = "_";
mem[41] = "_";
mem[42] = "_";
mem[43] = " ";
mem[44] = " ";
mem[45] = " ";
mem[46] = "\015";
mem[47] = "\012";
mem[48] = " ";
mem[49] = " ";
mem[50] = " ";
mem[51] = " ";
mem[52] = " ";
mem[53] = " ";
mem[54] = " ";
mem[55] = " ";
mem[56] = " ";
mem[57] = " ";
mem[58] = "d";
mem[59] = "e";
mem[60] = "l";
mem[61] = "a";
mem[62] = "y";
mem[63] = " ";
mem[64] = " ";
mem[65] = " ";
mem[66] = " ";
mem[67] = " ";
mem[68] = " ";
mem[69] = " ";
mem[70] = " ";
mem[71] = " ";
mem[72] = "|";
mem[73] = " ";
mem[74] = " ";
mem[75] = " ";
mem[76] = " ";
mem[77] = " ";
mem[78] = "p";
mem[79] = "u";
mem[80] = "l";
mem[81] = "s";
mem[82] = "e";
mem[83] = " ";
mem[84] = " ";
mem[85] = " ";
mem[86] = " ";
mem[87] = "|";
mem[88] = " ";
mem[89] = " ";
mem[90] = "\015";
mem[91] = "\012";
mem[92] = " ";
mem[93] = " ";
mem[94] = " ";
mem[95] = " ";
mem[96] = " ";
mem[97] = " ";
mem[98] = " ";
mem[99] = " ";
mem[100] = " ";
mem[101] = " ";
mem[102] = "w";
mem[103] = "i";
mem[104] = "d";
mem[105] = "t";
mem[106] = "h";
mem[107] = " ";
mem[108] = " ";
mem[109] = " ";
mem[110] = " ";
mem[111] = " ";
mem[112] = " ";
mem[113] = " ";
mem[114] = " ";
mem[115] = " ";
mem[116] = "|";
mem[117] = " ";
mem[118] = " ";
mem[119] = " ";
mem[120] = " ";
mem[121] = " ";
mem[122] = "w";
mem[123] = "i";
mem[124] = "d";
mem[125] = "t";
mem[126] = "h";
mem[127] = " ";
mem[128] = " ";
mem[129] = " ";
mem[130] = " ";
mem[131] = "|";
mem[132] = " ";
mem[133] = " ";
mem[134] = "\015";
mem[135] = "\012";
mem[136] = " ";
mem[137] = " ";
mem[138] = " ";
mem[139] = " ";
mem[140] = " ";
mem[141] = " ";
mem[142] = "";
mem[143] = "[";
mem[144] = "4";
mem[145] = "8";
mem[146] = ";";
mem[147] = "5";
mem[148] = ";";
mem[149] = "2";
mem[150] = "3";
mem[151] = "3";
mem[152] = "m";
mem[153] = " ";
mem[154] = " ";
mem[155] = "1";
mem[156] = "2";
mem[157] = "3";
mem[158] = "4";
mem[159] = "5";
mem[160] = "6";
mem[161] = "7";
mem[162] = "8";
mem[163] = " ";
mem[164] = " ";
mem[165] = "";
mem[166] = "[";
mem[167] = "m";
mem[168] = " ";
mem[169] = "n";
mem[170] = "s";
mem[171] = " ";
mem[172] = " ";
mem[173] = " ";
mem[174] = "|";
mem[175] = " ";
mem[176] = "";
mem[177] = "[";
mem[178] = "4";
mem[179] = "8";
mem[180] = ";";
mem[181] = "5";
mem[182] = ";";
mem[183] = "2";
mem[184] = "3";
mem[185] = "3";
mem[186] = "m";
mem[187] = " ";
mem[188] = " ";
mem[189] = "0";
mem[190] = "9";
mem[191] = "8";
mem[192] = "7";
mem[193] = "6";
mem[194] = "5";
mem[195] = "4";
mem[196] = "3";
mem[197] = " ";
mem[198] = " ";
mem[199] = "";
mem[200] = "[";
mem[201] = "m";
mem[202] = " ";
mem[203] = "|";
mem[204] = "n";
mem[205] = "s";
mem[206] = " ";
mem[207] = " ";
mem[208] = "\015";
mem[209] = "\012";
mem[210] = "_";
mem[211] = "_";
mem[212] = "_";
mem[213] = "_";
mem[214] = "_";
mem[215] = "_";
mem[216] = "_";
mem[217] = "_";
mem[218] = "_";
mem[219] = "_";
mem[220] = "_";
mem[221] = "_";
mem[222] = "_";
mem[223] = "_";
mem[224] = "_";
mem[225] = "_";
mem[226] = "_";
mem[227] = "_";
mem[228] = "_";
mem[229] = "_";
mem[230] = "_";
mem[231] = "_";
mem[232] = "_";
mem[233] = "_";
mem[234] = "|";
mem[235] = " ";
mem[236] = " ";
mem[237] = " ";
mem[238] = " ";
mem[239] = " ";
mem[240] = " ";
mem[241] = " ";
mem[242] = " ";
mem[243] = " ";
mem[244] = " ";
mem[245] = " ";
mem[246] = " ";
mem[247] = " ";
mem[248] = " ";
mem[249] = "|";
mem[250] = "_";
mem[251] = "_";
mem[252] = "\015";
mem[253] = "\012";
mem[254] = " ";
mem[255] = " ";
mem[256] = " ";
mem[257] = " ";
mem[258] = " ";
mem[259] = " ";
mem[260] = " ";
mem[261] = " ";
mem[262] = " ";
mem[263] = " ";
mem[264] = " ";
mem[265] = " ";
mem[266] = " ";
mem[267] = " ";
mem[268] = " ";
mem[269] = " ";
mem[270] = " ";
mem[271] = " ";
mem[272] = " ";
mem[273] = " ";
mem[274] = " ";
mem[275] = " ";
mem[276] = " ";
mem[277] = " ";
mem[278] = " ";
mem[279] = " ";
mem[280] = " ";
mem[281] = " ";
mem[282] = " ";
mem[283] = " ";
mem[284] = " ";
mem[285] = " ";
mem[286] = " ";
mem[287] = " ";
mem[288] = " ";
mem[289] = " ";
mem[290] = " ";
mem[291] = " ";
mem[292] = " ";
mem[293] = " ";
mem[294] = " ";
mem[295] = " ";
mem[296] = "\015";
mem[297] = "\012";
mem[298] = " ";
mem[299] = " ";
mem[300] = "t";
mem[301] = "a";
mem[302] = "b";
mem[303] = "=";
mem[304] = "f";
mem[305] = "i";
mem[306] = "e";
mem[307] = "l";
mem[308] = "d";
mem[309] = " ";
mem[310] = "s";
mem[311] = "p";
mem[312] = "a";
mem[313] = "c";
mem[314] = "e";
mem[315] = "=";
mem[316] = "r";
mem[317] = "e";
mem[318] = "d";
mem[319] = "r";
mem[320] = "a";
mem[321] = "w";
mem[322] = " ";
mem[323] = "e";
mem[324] = "n";
mem[325] = "t";
mem[326] = "e";
mem[327] = "r";
mem[328] = "=";
mem[329] = "t";
mem[330] = "r";
mem[331] = "i";
mem[332] = "g";
mem[333] = "g";
mem[334] = "e";
mem[335] = "r";
mem[336] = " ";
mem[337] = " ";
mem[338] = " ";
mem[339] = " ";
mem[340] = "\015";
mem[341] = "\012";
mem[342] = "";
mem[343] = "[";
mem[344] = "1";
mem[345] = ";";
mem[346] = "1";
mem[347] = "H";
