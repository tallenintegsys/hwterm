mem[0] = "K";
mem[1] = "N";
mem[2] = "O";
mem[3] = "W";
mem[4] = " ";
mem[5] = "A";
mem[6] = "L";
mem[7] = "L";
mem[8] = " ";
mem[9] = "M";
mem[10] = "E";
mem[11] = "N";
mem[12] = " ";
mem[13] = "B";
mem[14] = "Y";
mem[15] = " ";
mem[16] = "T";
mem[17] = "H";
mem[18] = "E";
mem[19] = "S";
mem[20] = "E";
mem[21] = " ";
mem[22] = "P";
mem[23] = "R";
mem[24] = "E";
mem[25] = "S";
mem[26] = "E";
mem[27] = "N";
mem[28] = "T";
mem[29] = "S";
mem[30] = ",";
mem[31] = " ";
mem[32] = "T";
mem[33] = "h";
mem[34] = "a";
mem[35] = "t";
mem[36] = " ";
mem[37] = "t";
mem[38] = "h";
mem[39] = "e";
mem[40] = " ";
mem[41] = "u";
mem[42] = "n";
mem[43] = "d";
mem[44] = "e";
mem[45] = "r";
mem[46] = "s";
mem[47] = "i";
mem[48] = "g";
mem[49] = "n";
mem[50] = "e";
mem[51] = "d";
mem[52] = ",";
mem[53] = " ";
mem[54] = "F";
mem[55] = "o";
mem[56] = "r";
mem[57] = " ";
mem[58] = "V";
mem[59] = "a";
mem[60] = "l";
mem[61] = "u";
mem[62] = "e";
mem[63] = " ";
mem[64] = "R";
mem[65] = "e";
mem[66] = "c";
mem[67] = "e";
mem[68] = "i";
mem[69] = "v";
mem[70] = "e";
mem[71] = "d";
mem[72] = ",";
mem[73] = " ";
mem[74] = "h";
mem[75] = "a";
mem[76] = "s";
mem[77] = " ";
mem[78] = "b";
mem[79] = "a";
mem[80] = "r";
mem[81] = "g";
mem[82] = "a";
mem[83] = "i";
mem[84] = "n";
mem[85] = "e";
mem[86] = "d";
mem[87] = ",";
mem[88] = " ";
mem[89] = "s";
mem[90] = "o";
mem[91] = "l";
mem[92] = "d";
mem[93] = ",";
mem[94] = " ";
mem[95] = "a";
mem[96] = "s";
mem[97] = "s";
mem[98] = "i";
mem[99] = "g";
mem[100] = "n";
mem[101] = "e";
mem[102] = "d";
mem[103] = " ";
mem[104] = "a";
mem[105] = "n";
mem[106] = "d";
mem[107] = " ";
mem[108] = "t";
mem[109] = "r";
mem[110] = "a";
mem[111] = "n";
mem[112] = "s";
mem[113] = "f";
mem[114] = "e";
mem[115] = "r";
mem[116] = "r";
mem[117] = "e";
mem[118] = "d";
mem[119] = " ";
mem[120] = "a";
mem[121] = "n";
mem[122] = "d";
mem[123] = " ";
mem[124] = "b";
mem[125] = "y";
mem[126] = " ";
mem[127] = "t";
mem[128] = "h";
mem[129] = "e";
mem[130] = "s";
mem[131] = "e";
mem[132] = " ";
mem[133] = "p";
mem[134] = "r";
mem[135] = "e";
mem[136] = "s";
mem[137] = "e";
mem[138] = "n";
mem[139] = "t";
mem[140] = "s";
mem[141] = " ";
mem[142] = "d";
mem[143] = "o";
mem[144] = "e";
mem[145] = "s";
mem[146] = " ";
mem[147] = "b";
mem[148] = "a";
mem[149] = "r";
mem[150] = "g";
mem[151] = "a";
mem[152] = "i";
mem[153] = "n";
mem[154] = ",";
mem[155] = " ";
mem[156] = "s";
mem[157] = "e";
mem[158] = "l";
mem[159] = "l";
mem[160] = ",";
mem[161] = " ";
mem[162] = "a";
mem[163] = "s";
mem[164] = "s";
mem[165] = "i";
mem[166] = "g";
mem[167] = "n";
mem[168] = " ";
mem[169] = "a";
mem[170] = "n";
mem[171] = "d";
mem[172] = " ";
mem[173] = "t";
mem[174] = "r";
mem[175] = "a";
mem[176] = "n";
mem[177] = "s";
mem[178] = "f";
mem[179] = "e";
mem[180] = "r";
mem[181] = " ";
mem[182] = "u";
mem[183] = "n";
mem[184] = "t";
mem[185] = "o";
mem[186] = " ";
mem[187] = "H";
mem[188] = "e";
mem[189] = "l";
mem[190] = "i";
mem[191] = "x";
mem[192] = " ";
mem[193] = "E";
mem[194] = "n";
mem[195] = "e";
mem[196] = "r";
mem[197] = "g";
mem[198] = "y";
mem[199] = " ";
mem[200] = "S";
mem[201] = "o";
mem[202] = "l";
mem[203] = "u";
mem[204] = "t";
mem[205] = "i";
mem[206] = "o";
mem[207] = "n";
mem[208] = "s";
mem[209] = " ";
mem[210] = "G";
mem[211] = "r";
mem[212] = "o";
mem[213] = "u";
mem[214] = "p";
mem[215] = ",";
mem[216] = " ";
mem[217] = "I";
mem[218] = "n";
mem[219] = "c";
mem[220] = ".";
mem[221] = ",";
mem[222] = " ";
mem[223] = "a";
mem[224] = " ";
mem[225] = "M";
mem[226] = "i";
mem[227] = "n";
mem[228] = "n";
mem[229] = "e";
mem[230] = "s";
mem[231] = "o";
mem[232] = "t";
mem[233] = "a";
mem[234] = " ";
mem[235] = "c";
mem[236] = "o";
mem[237] = "r";
mem[238] = "p";
mem[239] = "o";
mem[240] = "r";
mem[241] = "a";
mem[242] = "t";
mem[243] = "i";
mem[244] = "o";
mem[245] = "n";
mem[246] = " ";
mem[247] = "(";
mem[248] = "t";
mem[249] = "h";
mem[250] = "e";
mem[251] = " ";
mem[252] = "“";
mem[253] = "C";
mem[254] = "o";
mem[255] = "m";
mem[256] = "p";
mem[257] = "a";
mem[258] = "n";
mem[259] = "y";
mem[260] = "”";
mem[261] = ")";
mem[262] = ",";
mem[263] = " ";
mem[264] = "t";
mem[265] = "h";
mem[266] = "e";
mem[267] = " ";
mem[268] = "S";
mem[269] = "h";
mem[270] = "a";
mem[271] = "r";
mem[272] = "e";
mem[273] = "s";
mem[274] = " ";
mem[275] = "t";
mem[276] = "r";
mem[277] = "a";
mem[278] = "n";
mem[279] = "s";
mem[280] = "f";
mem[281] = "e";
mem[282] = "r";
mem[283] = "r";
mem[284] = "e";
mem[285] = "d";
mem[286] = " ";
mem[287] = "p";
mem[288] = "u";
mem[289] = "r";
mem[290] = "s";
mem[291] = "u";
mem[292] = "a";
mem[293] = "n";
mem[294] = "t";
mem[295] = " ";
mem[296] = "t";
mem[297] = "o";
mem[298] = " ";
mem[299] = "t";
mem[300] = "h";
mem[301] = "e";
mem[302] = " ";
mem[303] = "R";
mem[304] = "e";
mem[305] = "s";
mem[306] = "t";
mem[307] = "r";
mem[308] = "i";
mem[309] = "c";
mem[310] = "t";
mem[311] = "e";
mem[312] = "d";
mem[313] = " ";
mem[314] = "S";
mem[315] = "t";
mem[316] = "o";
mem[317] = "c";
mem[318] = "k";
mem[319] = " ";
mem[320] = "A";
mem[321] = "w";
mem[322] = "a";
mem[323] = "r";
mem[324] = "d";
mem[325] = " ";
mem[326] = "A";
mem[327] = "g";
mem[328] = "r";
mem[329] = "e";
mem[330] = "e";
mem[331] = "m";
mem[332] = "e";
mem[333] = "n";
mem[334] = "t";
mem[335] = " ";
mem[336] = "d";
mem[337] = "a";
mem[338] = "t";
mem[339] = "e";
mem[340] = "d";
mem[341] = " ";
mem[342] = "e";
mem[343] = "f";
mem[344] = "f";
mem[345] = "e";
mem[346] = "c";
mem[347] = "t";
mem[348] = "i";
mem[349] = "v";
mem[350] = "e";
mem[351] = " ";
mem[352] = "D";
mem[353] = "a";
mem[354] = "t";
mem[355] = "e";
mem[356] = ",";
mem[357] = " ";
mem[358] = "b";
mem[359] = "e";
mem[360] = "t";
mem[361] = "w";
mem[362] = "e";
mem[363] = "e";
mem[364] = "n";
mem[365] = " ";
mem[366] = "t";
mem[367] = "h";
mem[368] = "e";
mem[369] = " ";
mem[370] = "C";
mem[371] = "o";
mem[372] = "m";
mem[373] = "p";
mem[374] = "a";
mem[375] = "n";
mem[376] = "y";
mem[377] = " ";
mem[378] = "a";
mem[379] = "n";
mem[380] = "d";
mem[381] = " ";
mem[382] = "t";
mem[383] = "h";
mem[384] = "e";
mem[385] = " ";
mem[386] = "u";
mem[387] = "n";
mem[388] = "d";
mem[389] = "e";
mem[390] = "r";
mem[391] = "s";
mem[392] = "i";
mem[393] = "g";
mem[394] = "n";
mem[395] = "e";
mem[396] = "d";
mem[397] = ";";
mem[398] = " ";
mem[399] = "a";
mem[400] = "n";
mem[401] = "d";
mem[402] = " ";
mem[403] = "s";
mem[404] = "u";
mem[405] = "b";
mem[406] = "j";
mem[407] = "e";
mem[408] = "c";
mem[409] = "t";
mem[410] = " ";
mem[411] = "t";
mem[412] = "o";
mem[413] = " ";
mem[414] = "a";
mem[415] = "n";
mem[416] = "d";
mem[417] = " ";
mem[418] = "i";
mem[419] = "n";
mem[420] = " ";
mem[421] = "a";
mem[422] = "c";
mem[423] = "c";
mem[424] = "o";
mem[425] = "r";
mem[426] = "d";
mem[427] = "a";
mem[428] = "n";
mem[429] = "c";
mem[430] = "e";
mem[431] = " ";
mem[432] = "w";
mem[433] = "i";
mem[434] = "t";
mem[435] = "h";
mem[436] = " ";
mem[437] = "s";
mem[438] = "u";
mem[439] = "c";
mem[440] = "h";
mem[441] = " ";
mem[442] = "R";
mem[443] = "e";
mem[444] = "s";
mem[445] = "t";
mem[446] = "r";
mem[447] = "i";
mem[448] = "c";
mem[449] = "t";
mem[450] = "e";
mem[451] = "d";
mem[452] = " ";
mem[453] = "S";
mem[454] = "t";
mem[455] = "o";
mem[456] = "c";
mem[457] = "k";
mem[458] = " ";
mem[459] = "A";
mem[460] = "w";
mem[461] = "a";
mem[462] = "r";
mem[463] = "d";
mem[464] = " ";
mem[465] = "A";
mem[466] = "g";
mem[467] = "r";
mem[468] = "e";
mem[469] = "e";
mem[470] = "m";
mem[471] = "e";
mem[472] = "n";
mem[473] = "t";
mem[474] = " ";
mem[475] = "t";
mem[476] = "h";
mem[477] = "e";
mem[478] = " ";
mem[479] = "u";
mem[480] = "n";
mem[481] = "d";
mem[482] = "e";
mem[483] = "r";
mem[484] = "s";
mem[485] = "i";
mem[486] = "g";
mem[487] = "n";
mem[488] = "e";
mem[489] = "d";
mem[490] = " ";
mem[491] = "d";
mem[492] = "o";
mem[493] = "e";
mem[494] = "s";
mem[495] = " ";
mem[496] = "h";
mem[497] = "e";
mem[498] = "r";
mem[499] = "e";
mem[500] = "b";
mem[501] = "y";
mem[502] = " ";
mem[503] = "c";
mem[504] = "o";
mem[505] = "n";
mem[506] = "s";
mem[507] = "t";
mem[508] = "i";
mem[509] = "t";
mem[510] = "u";
mem[511] = "t";
mem[512] = "e";
mem[513] = " ";
mem[514] = "a";
mem[515] = "n";
mem[516] = "d";
mem[517] = " ";
mem[518] = "a";
mem[519] = "p";
mem[520] = "p";
mem[521] = "o";
mem[522] = "i";
mem[523] = "n";
mem[524] = "t";
mem[525] = " ";
mem[526] = "t";
mem[527] = "h";
mem[528] = "e";
mem[529] = " ";
mem[530] = "S";
mem[531] = "e";
mem[532] = "c";
mem[533] = "r";
mem[534] = "e";
mem[535] = "t";
mem[536] = "a";
mem[537] = "r";
mem[538] = "y";
mem[539] = " ";
mem[540] = "o";
mem[541] = "f";
mem[542] = " ";
mem[543] = "t";
mem[544] = "h";
mem[545] = "e";
mem[546] = " ";
mem[547] = "C";
mem[548] = "o";
mem[549] = "m";
mem[550] = "p";
mem[551] = "a";
mem[552] = "n";
mem[553] = "y";
mem[554] = " ";
mem[555] = "t";
mem[556] = "h";
mem[557] = "e";
mem[558] = " ";
mem[559] = "u";
mem[560] = "n";
mem[561] = "d";
mem[562] = "e";
mem[563] = "r";
mem[564] = "s";
mem[565] = "i";
mem[566] = "g";
mem[567] = "n";
mem[568] = "e";
mem[569] = "d";
mem[570] = "’";
mem[571] = "s";
mem[572] = " ";
mem[573] = "t";
mem[574] = "r";
mem[575] = "u";
mem[576] = "e";
mem[577] = " ";
mem[578] = "a";
mem[579] = "n";
mem[580] = "d";
mem[581] = " ";
mem[582] = "l";
mem[583] = "a";
mem[584] = "w";
mem[585] = "f";
mem[586] = "u";
mem[587] = "l";
mem[588] = " ";
mem[589] = "a";
mem[590] = "t";
mem[591] = "t";
mem[592] = "o";
mem[593] = "r";
mem[594] = "n";
mem[595] = "e";
mem[596] = "y";
mem[597] = ",";
mem[598] = " ";
mem[599] = "I";
mem[600] = "R";
mem[601] = "R";
mem[602] = "E";
mem[603] = "V";
mem[604] = "O";
mem[605] = "C";
mem[606] = "A";
mem[607] = "B";
mem[608] = "L";
mem[609] = "Y";
mem[610] = ",";
mem[611] = " ";
mem[612] = "t";
mem[613] = "o";
mem[614] = " ";
mem[615] = "s";
mem[616] = "e";
mem[617] = "l";
mem[618] = "l";
mem[619] = " ";
mem[620] = "a";
mem[621] = "s";
mem[622] = "s";
mem[623] = "i";
mem[624] = "g";
mem[625] = "n";
mem[626] = ",";
mem[627] = " ";
mem[628] = "t";
mem[629] = "r";
mem[630] = "a";
mem[631] = "n";
mem[632] = "s";
mem[633] = "f";
mem[634] = "e";
mem[635] = "r";
mem[636] = ",";
mem[637] = " ";
mem[638] = "h";
mem[639] = "y";
mem[640] = "p";
mem[641] = "o";
mem[642] = "t";
mem[643] = "h";
mem[644] = "e";
mem[645] = "c";
mem[646] = "a";
mem[647] = "t";
mem[648] = "e";
mem[649] = ",";
mem[650] = " ";
mem[651] = "p";
mem[652] = "l";
mem[653] = "e";
mem[654] = "d";
mem[655] = "g";
mem[656] = "e";
mem[657] = " ";
mem[658] = "a";
mem[659] = "n";
mem[660] = "d";
mem[661] = " ";
mem[662] = "m";
mem[663] = "a";
mem[664] = "k";
mem[665] = "e";
mem[666] = " ";
mem[667] = "o";
mem[668] = "v";
mem[669] = "e";
mem[670] = "r";
mem[671] = " ";
mem[672] = "a";
mem[673] = "l";
mem[674] = "l";
mem[675] = " ";
mem[676] = "o";
mem[677] = "r";
mem[678] = " ";
mem[679] = "a";
mem[680] = "n";
mem[681] = "y";
mem[682] = " ";
mem[683] = "p";
mem[684] = "a";
mem[685] = "r";
mem[686] = "t";
mem[687] = " ";
mem[688] = "o";
mem[689] = "f";
mem[690] = " ";
mem[691] = "s";
mem[692] = "u";
mem[693] = "c";
mem[694] = "h";
mem[695] = " ";
mem[696] = "S";
mem[697] = "h";
mem[698] = "a";
mem[699] = "r";
mem[700] = "e";
mem[701] = "s";
mem[702] = " ";
mem[703] = "a";
mem[704] = "n";
mem[705] = "d";
mem[706] = " ";
mem[707] = "f";
mem[708] = "o";
mem[709] = "r";
mem[710] = " ";
mem[711] = "t";
mem[712] = "h";
mem[713] = "a";
mem[714] = "t";
mem[715] = " ";
mem[716] = "p";
mem[717] = "u";
mem[718] = "r";
mem[719] = "p";
mem[720] = "o";
mem[721] = "s";
mem[722] = "e";
mem[723] = " ";
mem[724] = "t";
mem[725] = "o";
mem[726] = " ";
mem[727] = "m";
mem[728] = "a";
mem[729] = "k";
mem[730] = "e";
mem[731] = " ";
mem[732] = "a";
mem[733] = "n";
mem[734] = "d";
mem[735] = " ";
mem[736] = "e";
mem[737] = "x";
mem[738] = "e";
mem[739] = "c";
mem[740] = "u";
mem[741] = "t";
mem[742] = "e";
mem[743] = " ";
mem[744] = "a";
mem[745] = "l";
mem[746] = "l";
mem[747] = " ";
mem[748] = "n";
mem[749] = "e";
mem[750] = "c";
mem[751] = "e";
mem[752] = "s";
mem[753] = "s";
mem[754] = "a";
mem[755] = "r";
mem[756] = "y";
mem[757] = " ";
mem[758] = "a";
mem[759] = "c";
mem[760] = "t";
mem[761] = "s";
mem[762] = " ";
mem[763] = "o";
mem[764] = "f";
mem[765] = " ";
mem[766] = "a";
mem[767] = "s";
mem[768] = "s";
mem[769] = "i";
mem[770] = "g";
mem[771] = "n";
mem[772] = "m";
mem[773] = "e";
mem[774] = "n";
mem[775] = "t";
mem[776] = " ";
mem[777] = "a";
mem[778] = "n";
mem[779] = "d";
mem[780] = " ";
mem[781] = "t";
mem[782] = "r";
mem[783] = "a";
mem[784] = "n";
mem[785] = "s";
mem[786] = "f";
mem[787] = "e";
mem[788] = "r";
mem[789] = " ";
mem[790] = "t";
mem[791] = "h";
mem[792] = "e";
mem[793] = "r";
mem[794] = "e";
mem[795] = "o";
mem[796] = "f";
mem[797] = ",";
mem[798] = " ";
mem[799] = "a";
mem[800] = "n";
mem[801] = "d";
mem[802] = " ";
mem[803] = "t";
mem[804] = "o";
mem[805] = " ";
mem[806] = "s";
mem[807] = "u";
mem[808] = "b";
mem[809] = "s";
mem[810] = "t";
mem[811] = "i";
mem[812] = "t";
mem[813] = "u";
mem[814] = "t";
mem[815] = "e";
mem[816] = " ";
mem[817] = "o";
mem[818] = "n";
mem[819] = "e";
mem[820] = " ";
mem[821] = "o";
mem[822] = "r";
mem[823] = " ";
mem[824] = "m";
mem[825] = "o";
mem[826] = "r";
mem[827] = "e";
mem[828] = " ";
mem[829] = "p";
mem[830] = "e";
mem[831] = "r";
mem[832] = "s";
mem[833] = "o";
mem[834] = "n";
mem[835] = "s";
mem[836] = " ";
mem[837] = "w";
mem[838] = "i";
mem[839] = "t";
mem[840] = "h";
mem[841] = " ";
mem[842] = "l";
mem[843] = "i";
mem[844] = "k";
mem[845] = "e";
mem[846] = " ";
mem[847] = "f";
mem[848] = "u";
mem[849] = "l";
mem[850] = "l";
mem[851] = " ";
mem[852] = "p";
mem[853] = "o";
mem[854] = "w";
mem[855] = "e";
mem[856] = "r";
mem[857] = ",";
mem[858] = " ";
mem[859] = "h";
mem[860] = "e";
mem[861] = "r";
mem[862] = "e";
mem[863] = "b";
mem[864] = "y";
mem[865] = " ";
mem[866] = "r";
mem[867] = "a";
mem[868] = "t";
mem[869] = "i";
mem[870] = "f";
mem[871] = "y";
mem[872] = "i";
mem[873] = "n";
mem[874] = "g";
mem[875] = " ";
mem[876] = "a";
mem[877] = "n";
mem[878] = "d";
mem[879] = " ";
mem[880] = "c";
mem[881] = "o";
mem[882] = "n";
mem[883] = "f";
mem[884] = "i";
mem[885] = "r";
mem[886] = "m";
mem[887] = "i";
mem[888] = "n";
mem[889] = "g";
mem[890] = " ";
mem[891] = "a";
mem[892] = "l";
mem[893] = "l";
mem[894] = " ";
mem[895] = "t";
mem[896] = "h";
mem[897] = "a";
mem[898] = "t";
mem[899] = " ";
mem[900] = "s";
mem[901] = "a";
mem[902] = "i";
mem[903] = "d";
mem[904] = " ";
mem[905] = "a";
mem[906] = "t";
mem[907] = "t";
mem[908] = "o";
mem[909] = "r";
mem[910] = "n";
mem[911] = "e";
mem[912] = "y";
mem[913] = " ";
mem[914] = "o";
mem[915] = "r";
mem[916] = " ";
mem[917] = "h";
mem[918] = "i";
mem[919] = "s";
mem[920] = " ";
mem[921] = "s";
mem[922] = "u";
mem[923] = "b";
mem[924] = "s";
mem[925] = "t";
mem[926] = "i";
mem[927] = "t";
mem[928] = "u";
mem[929] = "t";
mem[930] = "e";
mem[931] = "s";
mem[932] = " ";
mem[933] = "s";
mem[934] = "h";
mem[935] = "a";
mem[936] = "l";
mem[937] = "l";
mem[938] = " ";
mem[939] = "l";
mem[940] = "a";
mem[941] = "w";
mem[942] = "f";
mem[943] = "u";
mem[944] = "l";
mem[945] = "l";
mem[946] = "y";
mem[947] = " ";
mem[948] = "d";
mem[949] = "o";
mem[950] = " ";
mem[951] = "b";
mem[952] = "y";
mem[953] = " ";
mem[954] = "v";
mem[955] = "i";
mem[956] = "r";
mem[957] = "t";
mem[958] = "u";
mem[959] = "e";
mem[960] = " ";
mem[961] = "h";
mem[962] = "e";
mem[963] = "r";
mem[964] = "e";
mem[965] = "o";
mem[966] = "f";
mem[967] = ".";
mem[968] = "I";
mem[969] = "t";
mem[970] = " ";
mem[971] = "o";
mem[972] = "c";
mem[973] = "c";
mem[974] = "u";
mem[975] = "r";
mem[976] = "s";
mem[977] = " ";
mem[978] = "i";
mem[979] = "n";
mem[980] = " ";
mem[981] = "b";
mem[982] = "i";
mem[983] = "l";
mem[984] = "l";
mem[985] = "s";
mem[986] = " ";
mem[987] = "o";
mem[988] = "f";
mem[989] = " ";
mem[990] = "s";
mem[991] = "a";
mem[992] = "l";
mem[993] = "e";
mem[994] = ",";
mem[995] = " ";
mem[996] = "i";
mem[997] = "n";
mem[998] = "s";
mem[999] = "t";
mem[1000] = "r";
mem[1001] = "u";
mem[1002] = "m";
mem[1003] = "e";
mem[1004] = "n";
mem[1005] = "t";
mem[1006] = "s";
mem[1007] = " ";
mem[1008] = "o";
mem[1009] = "f";
mem[1010] = " ";
mem[1011] = "a";
mem[1012] = "s";
mem[1013] = "s";
mem[1014] = "i";
mem[1015] = "g";
mem[1016] = "n";
mem[1017] = "m";
mem[1018] = "e";
mem[1019] = "n";
mem[1020] = "t";
mem[1021] = ",";
mem[1022] = " ";
mem[1023] = "r";
